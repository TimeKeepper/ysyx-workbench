import "DPI-C" function int npc_trap (input int ra);

module sram(
    input clock,
    input reset,
    input [31:0] addr,
    input [31:0] w_data,
    input w_r,

    output [31:0] r_data,
    output valid
)



endmodule