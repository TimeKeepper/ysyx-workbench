module work(
    input clk,
    input rst,
    output [15:0] mem_store
);

    

endmodule